`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/22/2020 12:52:41 PM
// Design Name: 
// Module Name: reg_define
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


// $Id$
// This file was generated by regmaker.pl

module reg_define (
    output reg [1:0]  turn_on_signal, // start_sytolic_array 
    output reg [31:0] input_acc_size, // input_acc_size 

    input      [31:0] write_data,
    input      [15:0] addr,
    output     [31:0] read_data,
    input write,
    input read,
    input clk,
    input reset_l
     );

wire [15:0] addr_1;
wire [31:0] write_data_1;
reg  [31:0] read_data_1;
wire read_1, write_1;

assign addr_1       = addr;
assign write_data_1 = write_data;
assign write_1      = write;
assign read_1       = read;
assign read_data    = read_data_1;


// read data is available in the same cycle as when addr is applied
// write data is available 1 cycle after addr is applied

always @(posedge clk or negedge reset_l) begin
    if (!reset_l) begin
        turn_on_signal <= 2'h0; // turn on the hese encoder and comparator
        input_acc_size <= 32'h00000000; // input_acc_size 
     end
    else begin

      if (write_1) begin
        case(addr_1[15:0])
            16'h0000: begin  // start_sytolic_array
                turn_on_signal[1:0] <= write_data_1[1:0];
            end
            16'h0008: begin  // input_acc_size
                input_acc_size[31:0] <= write_data_1[31:0];
            end

        endcase
    end
  end
end
// Reads...
       always @* begin
           case(addr_1[15:0])
              16'h0004: begin // sytolic_array_idle
                read_data_1 = {30'h00000000,turn_on_signal[1:0]};
              end
              16'h0008: begin // input_acc_size
                read_data_1 = {input_acc_size[31:0]};
              end

              default: read_data_1 = {16'hdead,addr_1[15:0]};
          endcase
      end

endmodule

